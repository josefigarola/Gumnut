module Stack(
	//de a egg globales
	input logic clk,
	input logic cen,
	input logic rst,
	input logic pop_i,
	input logic push_i,
	input logic [11:0]pc_i, //viene de progcounter
	//output
	output logic [11:0]spc_o
	);
	
endmodule 